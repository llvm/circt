// This module is used in the library locations test.
// Empty `RUN` line such that it does not get picked up by lit.
// RUN:

module library_module;
endmodule
