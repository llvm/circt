module ExtResource(); endmodule
