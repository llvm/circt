module Bar();
endmodule
