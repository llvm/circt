module ifdef(output out);
   assign out = 1'b1;
endmodule
