// This file is included from `preprocess.sv`. Empty `RUN` line such that it
// does not get picked up by lit.
// RUN:

localparam Z = 9001;
