// REQUIRES: verilator
// RUN: verilator --cc --top-module basics -Wall -Wpedantic %s

module basics ();

endmodule
